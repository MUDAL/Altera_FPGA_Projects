library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

-- Package that contains constants and function(s) that ....
-- are relevant to the project.

package pkg is
   function log_base2(param: integer) return integer;
   -- Memory Initialization File (MIF) parameters
   constant MIF_LEN:       integer := 24;
   constant GAME_MENU_MIF: string(1 to MIF_LEN) := "../src/mif/game_menu.mif";
   constant GAME_OVER_MIF: string(1 to MIF_LEN) := "../src/mif/game_over.mif";
   ------------------------------------------------------------------
   -- Ball Directions
   constant DIR_UR: std_logic_vector(2 downto 0) := "000"; -- Up + Right
   constant DIR_R:  std_logic_vector(2 downto 0) := "001"; -- Right
   constant DIR_DR: std_logic_vector(2 downto 0) := "010"; -- Down + Right
   constant DIR_DL: std_logic_vector(2 downto 0) := "011"; -- Down + Left
   constant DIR_L:  std_logic_vector(2 downto 0) := "100"; -- Left
   constant DIR_UL: std_logic_vector(2 downto 0) := "101"; -- Up + Left
   ------------------------------------------------------------------
   -- Number of rows and columns for the fonts [Powers of 2 are recommended]
   constant COLS: integer := 8;
   constant ROWS: integer := 8;  
   ------------------------------------------------------------------
   -- Font Type Declaration
   type font_t is array(0 to ROWS - 1) of std_logic_vector(0 to COLS - 1);
   ------------------------------------------------------------------
   constant FONT_0: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "01000010",
                               4 => "01000010",
                               5 => "01000010",
                               6 => "01111110",
                               7 => "00000000");   
   ------------------------------------------------------------------  
   constant FONT_1: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "00000010",
                               3 => "00000010",
                               4 => "00000010",
                               5 => "00000010",
                               6 => "00000010",
                               7 => "00000000");
   ------------------------------------------------------------------    
   constant FONT_2: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "00000010",
                               4 => "01111110",
                               5 => "01000000",
                               6 => "01111110",
                               7 => "00000000");
   ------------------------------------------------------------------    
   constant FONT_3: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "00000010",
                               4 => "01111110",
                               5 => "00000010",
                               6 => "01111110",
                               7 => "00000000");
   ------------------------------------------------------------------   
   constant FONT_4: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01000010",
                               3 => "01000010",
                               4 => "01111110",
                               5 => "00000010",
                               6 => "00000010",
                               7 => "00000000");
   ------------------------------------------------------------------                               
   constant FONT_5: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "01000000",
                               4 => "01111110",
                               5 => "00000010",
                               6 => "01111110",
                               7 => "00000000");
   ------------------------------------------------------------------
   constant FONT_6: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "01000000",
                               4 => "01111110",
                               5 => "01000010",
                               6 => "01111110",
                               7 => "00000000");   
   ------------------------------------------------------------------                            
   constant FONT_7: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "00000010",
                               4 => "00000010",
                               5 => "00000010",
                               6 => "00000010",
                               7 => "00000000");
   ------------------------------------------------------------------
   constant FONT_8: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "01000010",
                               4 => "01111110",
                               5 => "01000010",
                               6 => "01111110",
                               7 => "00000000");
   ------------------------------------------------------------------                            
   constant FONT_9: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "01111110",
                               3 => "01000010",
                               4 => "01111110",
                               5 => "00000010",
                               6 => "01111110",
                               7 => "00000000");                                  
   ------------------------------------------------------------------                            
   constant F_NULL: font_t := (0 => "00000000",
                               1 => "00000000",
                               2 => "00000000",
                               3 => "00000000",
                               4 => "00000000",
                               5 => "00000000",
                               6 => "00000000",
                               7 => "00000000");                               
   ------------------------------------------------------------------
   constant ROM_DEPTH:      integer := 16;
   constant DIG_ADDR_WIDTH: integer := 4; -- Address width for digits in ROM
   ------------------------------------------------------------------
   -- Font ROM
   type rom_t is array(0 to ROM_DEPTH - 1) of font_t;   
   constant ROM: rom_t := (0 => FONT_0,
                           1 => FONT_1,
                           2 => FONT_2,
                           3 => FONT_3,
                           4 => FONT_4,
                           5 => FONT_5,
                           6 => FONT_6,
                           7 => FONT_7,
                           8 => FONT_8,
                           9 => FONT_9,
                           others => F_NULL);
   ------------------------------------------------------------------                           
end package pkg;

---------------------------------------------------------------------
--                         PACKAGE BODY
---------------------------------------------------------------------

package body pkg is
   ------------------------------------------------------------------
   function log_base2(param: integer) return integer is
   begin
      return integer(ceil(log2(real(param))));
   end function log_base2;
   ------------------------------------------------------------------
end package body pkg;